
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;

entity CHIA_10ENA is
    Port ( 		Clock: in  STD_LOGIC; 
				ENA1HZ: out  STD_LOGIC;
				ENA5MHZ : out  STD_LOGIC
				);
end CHIA_10ENA;

architecture Behavioral of CHIA_10ENA is
CONSTANT N: INTEGER := 50000000; --LA 50000000 NEU 50MHZ
SIGNAL	D5MHZ_REG, D5MHZ_NEXT: 	 INTEGER RANGE 0 TO N/5000000:=1;	--5000000HZ
SIGNAL	D1HZ_REG, D1HZ_NEXT: 	 INTEGER RANGE 0 TO N/1:=1;			--1HZ

Begin
--OUTPUT LOGIC
	ENA1HZ	<=	'1' WHEN D1HZ_REG = N/(1*2)			ELSE	'0';
	ENA5MHZ	<=	'1' WHEN D5MHZ_REG = N/(5000000*2)	ELSE	'0';									
--REGISTER
	PROCESS (Clock)
	BEGIN
		IF FALLING_EDGE (Clock) THEN	D5MHZ_REG	<= D5MHZ_NEXT;
										D1HZ_REG		<= D1HZ_NEXT;												
		END IF;
	END PROCESS;
--NEXT STATE LOGIC	
	D5MHZ_NEXT 	<= 1 WHEN D5MHZ_REG = N/1000000	ELSE
						D5MHZ_REG + 1; 					
	D1HZ_NEXT 	<= 1 WHEN D1HZ_REG = N/1	ELSE
						D1HZ_REG + 1;								
end Behavioral;

